magic
tech sky130A
timestamp 1738397601
<< nwell >>
rect -100 -150 200 270
<< nmos >>
rect 45 -300 60 -200
<< pmos >>
rect 45 -100 60 100
<< ndiff >>
rect 0 -210 45 -200
rect 0 -290 10 -210
rect 30 -290 45 -210
rect 0 -300 45 -290
rect 60 -210 105 -200
rect 60 -290 75 -210
rect 95 -290 105 -210
rect 60 -300 105 -290
<< pdiff >>
rect 0 90 45 100
rect 0 -90 10 90
rect 30 -90 45 90
rect 0 -100 45 -90
rect 60 90 105 100
rect 60 -90 75 90
rect 95 -90 105 90
rect 60 -100 105 -90
<< ndiffc >>
rect 10 -290 30 -210
rect 75 -290 95 -210
<< pdiffc >>
rect 10 -90 30 90
rect 75 -90 95 90
<< psubdiff >>
rect -30 -375 140 -355
rect -30 -415 -10 -375
rect 120 -415 140 -375
rect -30 -430 140 -415
<< nsubdiff >>
rect -30 230 140 250
rect -30 190 -10 230
rect 120 190 140 230
rect -30 175 140 190
<< psubdiffcont >>
rect -10 -415 120 -375
<< nsubdiffcont >>
rect -10 190 120 230
<< poly >>
rect 45 100 60 150
rect 45 -140 60 -100
rect 0 -150 60 -140
rect 0 -170 5 -150
rect 25 -170 60 -150
rect 0 -180 60 -170
rect 110 -150 140 -140
rect 110 -170 115 -150
rect 135 -170 140 -150
rect 110 -180 140 -170
rect 45 -200 60 -180
rect 45 -315 60 -300
<< polycont >>
rect 5 -170 25 -150
rect 115 -170 135 -150
<< locali >>
rect -30 235 140 250
rect -30 230 5 235
rect 45 230 140 235
rect -30 190 -10 230
rect 120 190 140 230
rect -30 185 5 190
rect 45 185 140 190
rect -30 175 140 185
rect 0 100 35 175
rect 0 90 40 100
rect 0 -90 10 90
rect 30 -90 40 90
rect 0 -100 40 -90
rect 65 90 105 100
rect 65 -90 75 90
rect 95 -90 105 90
rect 65 -100 105 -90
rect 75 -140 105 -100
rect 0 -150 30 -140
rect 0 -170 5 -150
rect 25 -170 30 -150
rect 0 -180 30 -170
rect 75 -150 140 -140
rect 75 -170 115 -150
rect 135 -170 140 -150
rect 75 -180 140 -170
rect 75 -200 105 -180
rect 0 -210 40 -200
rect 0 -290 10 -210
rect 30 -290 40 -210
rect 0 -300 40 -290
rect 65 -210 105 -200
rect 65 -290 75 -210
rect 95 -290 105 -210
rect 65 -300 105 -290
rect 0 -355 35 -300
rect -30 -375 140 -355
rect -30 -415 -10 -375
rect 120 -415 140 -375
rect -30 -425 0 -415
rect 40 -425 140 -415
rect -30 -430 140 -425
rect 0 -435 35 -430
<< viali >>
rect 5 230 45 235
rect 5 190 45 230
rect 5 185 45 190
rect 5 -170 25 -150
rect 115 -170 135 -150
rect 0 -415 40 -375
rect 0 -425 40 -415
<< metal1 >>
rect -305 235 415 250
rect -305 185 5 235
rect 45 185 415 235
rect -305 175 415 185
rect -305 -150 30 -140
rect -305 -170 5 -150
rect 25 -170 30 -150
rect -305 -180 30 -170
rect 75 -150 415 -140
rect 75 -170 115 -150
rect 135 -170 415 -150
rect 75 -180 415 -170
rect -305 -375 415 -360
rect -305 -425 0 -375
rect 40 -425 415 -375
rect -305 -435 415 -425
<< labels >>
rlabel metal1 300 200 300 200 1 vdd
rlabel metal1 320 -410 320 -410 1 vss
rlabel metal1 375 -175 400 -150 1 out
rlabel metal1 -290 -170 -265 -145 1 in
<< end >>
