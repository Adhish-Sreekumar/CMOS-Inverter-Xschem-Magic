* SPICE3 file created from /home/vboxuser/Desktop/first_test/magic_tests/inverter_scratch.ext - technology: sky130A

X0 out in vss vss sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X1 out in vdd vdd sky130_fd_pr__pfet_01v8 ad=0.9 pd=4.9 as=0.9 ps=4.9 w=2 l=0.15
C0 vdd vss 2.20771f **FLOATING
